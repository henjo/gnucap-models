flux shuttle shift register
r1 1 2 100
r2 2 0 .4
r3 3 0 .4
r4 4 0 .4
r5 5 0 .4
r6 6 0 .4
r7 7 0 .4
r8 8 0 .4
r9 9 0 .4
r10 10 11 100
r20 20 21 100
r30 30 31 100

l1 2 3 3p
l2 3 4 3p
l3 4 5 3p
l4 5 6 3p
l5 6 7 3p
l6 7 8 3p
l7 8 9 3p

l10 11 12 3p
l11 12 13 3p
l12 13 0  3p
l20 21 22 3p
l21 22 0  3p
l30 31 32 3p
l31 32 0  3p

k1 l10 l1 .99
k2 l11 l4 .99
k3 l12 l7 .99
k4 l20 l2 .99
k5 l21 l5 .99
k6 l30 l3 .99
k7 l31 l6 .99

b1 2 0 100 jj1
b2 3 0 101 jj1
b3 4 0 102 jj1
b4 5 0 103 jj1
b5 6 0 104 jj1
b6 7 0 105 jj1
b7 8 0 106 jj1
b8 9 0 107 jj1

* couple phi2 into last junction to clear
rxx 9 20 140

*v1 10 0 pulse(0 120m  25p 10p 10p 10p 120p)
*v2 20 0 pulse(0 120m  65p 10p 10p 10p 120p)
*v3 30 0 pulse(0 120m 105p 10p 10p 10p 120p)
*v4 1 0 pulse(0 40m 25p 10p 10p)

v1 10 0 spulse(0 120m 120p 25p)
v2 20 0 spulse(0 120m 120p 65p)
v3 30 0 spulse(0 120m 120p 105p)
*v4 1 0 pulse(0 40m 15p 10p 10p 60p)
v4 1 0 pulse(0 30m 70p 10p 10p 10p 360p)
*v5 200 0 pulse(0 30m 430p 10p 10p 10p)

*Nb 2500 A/cm2   area = 40 square microns
.model jj1 jj(rtype=1,cct=1,icon=10m,vg=2.8m,delv=0.08m,
+ icrit=1m,r0=30,rn=1.647059,cap=1.548944p)
.end
